* SPICE3 file created from nand.ext - technology: scmos
.include tsmc_cmos025
.option scale=0.12u

.model nfet NMOS
.model pfet PMOS

Vdd vdd 0 2.5V
VinA A gnd PULSE(2.5 0 0ns 10ns 10ns 20ns 40ns)
VinB B gnd PULSE(2.5 0 0ns 5ns 10ns 20ns 40ns)
CL Z gnd 1fF
.TRAN 1ns 100ns

M1000 vdd B Z vdd pfet w=8 l=2
+  ad=80 pd=52 as=48 ps=28
M1001 Z A vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_n2_n41# A gnd gnd nfet w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1003 Z B a_n2_n41# gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 B A 0.33fF
C1 Z B 0.07fF
C2 vdd A 0.10fF
C3 vdd Z 0.25fF
C4 vdd B 0.10fF
C5 gnd Z 0.02fF
C6 Z A 0.05fF
C7 gnd gnd 0.13fF
C8 Z gnd 0.37fF
C9 B gnd 0.72fF
C10 A gnd 0.75fF
C11 vdd gnd 0.71fF

* Delay measurements for NAND2 gate
.measure tran tp_nand_a TRIG V(A) VAL=0.3 FALL=1 TARG V(Z) VAL=0.3 RISE=1
.measure tran tp_nand_b TRIG V(B) VAL=2 FALL=1 TARG V(Z) VAL=2 RISE=1

* Simulation control commands
.control
run
print tp_nand_a
print tp_nand_b
.endc

.end

