* SPICE3 file created from nor.ext - technology: scmos

.include tsmc_cmos025
.option scale=0.12u

.model nfet NMOS
.model pfet PMOS

Vdd vdd 0 2.5V
VinA A gnd PULSE(0 2.5 0ns 10ns 10ns 20ns 40ns)
VinB B gnd PULSE(0 2.5 0ns 5ns 10ns 20ns 40ns)
CL Z gnd 1fF
.TRAN 1ns 100ns

* Delay measurements for NAND2 gate
.measure tran tp_nand_a TRIG V(A) VAL=0.3 FALL=1 TARG V(Z) VAL=0.3 RISE=1
.measure tran tp_nand_b TRIG V(B) VAL=2 FALL=1 TARG V(Z) VAL=2 RISE=1

* Simulation control commands
.control
run
print tp_nand_a
print tp_nand_b
.endc

M1000 Z B a_n2_34# vdd pfet w=8 l=2
+  ad=40 pd=26 as=48 ps=28
M1001 Z A gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=40 ps=36
M1002 a_n2_34# A vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1003 gnd B Z Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A B 0.33fF
C1 gnd Z 0.12fF
C2 vdd B 0.10fF
C3 B Z 0.12fF
C4 vdd A 0.10fF
C5 vdd Z 0.08fF
C6 gnd Gnd 0.16fF
C7 Z Gnd 0.41fF
C8 B Gnd 0.73fF
C9 A Gnd 0.76fF
C10 vdd Gnd 0.71fF

.end
